--- ini untuk top dari top 
